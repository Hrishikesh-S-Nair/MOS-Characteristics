*pMOS Transfer Characteristics
vdd 2 0 dc 1.5v
vd 3 0 dc 0v
vgs 1 0 dc 2v
m1 2 1 0 3 pmos1 w=180n l=90n
.model pmos1 pmos vt0=1.5v kp=200u
.dc vdd 0 1.5 0.01
.control
set color0=white
run
plot i(vd) ylabel 'Ids' xlabel 'Vds' title 'Output Characteristics'
.endc
.end